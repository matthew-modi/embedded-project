module camera_interface (
    input logic clk,
    input logic reset,
    input logic [7:0] d,
    input logic href,
    input logic vsync
);

endmodule